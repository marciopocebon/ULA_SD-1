module CPU(barramento, Tx,Ty,Tz,Tula, clock, a, b, saidaULA, saida)
    input wire clock;
    output [3:0] barramento;
    
endmodule